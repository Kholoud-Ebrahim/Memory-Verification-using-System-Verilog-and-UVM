package utils_pkg;
	parameter DATA_WIDTH = 32;
  parameter ADDR_WIDTH = 4;
endpackage:utils_pkg
